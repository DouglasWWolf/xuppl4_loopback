/*
================================================================================================
   Vers    Date     Who  Changes
 ------  ---------------------------------------------------------------------------------------
  1.0.1  04-Jun-24  DWW  Initial creation
  1.1.0  08-Jun-24  DWW  Added run-time configurability of RS-FEC and TX pre-emphasis
  1.2.0  15-Jun-24  DWW  Now controlling CMAC gt_txdiffctrl
  1.3.0  16-Jun-24  DWW  txpost and txdiff are now programmable
  1.3.1  30-Jun-24  DWW  Set SYSTEM_JITTER to 300ps to tighten up timing
  1.4.0  04-Jul-25  DWW  Integrated with the build system
================================================================================================
*/

localparam VERSION_MAJOR = 1;
localparam VERSION_MINOR = 4;
localparam VERSION_BUILD = 0;
localparam VERSION_RCAND = 0;

localparam RTL_TYPE      = 642024;
localparam RTL_SUBTYPE   = 0;


//================================================================================================
//    Date      Vers   Who  Changes
// -----------------------------------------------------------------------------------------------
// 04-Jun-2024  1.0.1  DWW  Initial creation
//================================================================================================
localparam VERSION_MAJOR = 1;
localparam VERSION_MINOR = 0;
localparam VERSION_BUILD = 1;
localparam VERSION_RCAND = 0;

localparam VERSION_DAY   = 4;
localparam VERSION_MONTH = 6;
localparam VERSION_YEAR  = 2024;

localparam RTL_TYPE      = 642024;
localparam RTL_SUBTYPE   = 0;
